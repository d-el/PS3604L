* D:\Radio\Devices\PS3608L\OrCad\CulerReg.sch

* Schematics Version 9.2
* Mon Aug 08 01:46:47 2016



** Analysis setup **
.tran 20ns 100ms


* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "CulerReg.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
