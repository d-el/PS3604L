** Profile: "SCHEMATIC1-Bias"  [ d:\radio\devices\ps3608l\orcad\str-schematic1-bias.sim ] 

** Creating circuit file "str-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:

*Analysis directives: 
.TRAN  0 1000ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\str-SCHEMATIC1.net" 


.END
