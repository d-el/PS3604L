* D:\Radio\Devices\PS3608L\OrCad\Rectifier.sch

* Schematics Version 9.2
* Thu Sep 29 20:54:08 2016



** Analysis setup **
.tran 20n 15m


* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Rectifier.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
