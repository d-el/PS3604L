** Profile: "SCHEMATIC1-timetrans"  [ D:\Radio\Devices\PS3604L\OrCad\outamp\outamp-SCHEMATIC1-timetrans.sim ] 

** Creating circuit file "outamp-SCHEMATIC1-timetrans.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\phil_bjt.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\anlg_dev.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\opamp.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\opamp.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\ediode.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\pwrmos.lib" 
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\diode.lib" 

*Analysis directives: 
.TRAN  0 2000us 0 1ms 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\outamp-SCHEMATIC1.net" 


.END
