** Profile: "SCHEMATIC1-timetrans1"  [ D:\Radio\Devices\PS3604L\OrCad\outamp\outamp-schematic1-timetrans1.sim ] 

** Creating circuit file "outamp-schematic1-timetrans1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\nom.lib" 
.inc "C:\ProgramFiles\Orcad\Capture\Library\PSpice\nom.lib" 

*Analysis directives: 
.TRAN  0 600000u 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\outamp-SCHEMATIC1.net" 


.END
