** Profile: "SCHEMATIC1-Trans"  [ D:\Radio\Devices\PS3604L\OrCad\rectifier\rectifier-schematic1-trans.sim ] 

** Creating circuit file "rectifier-schematic1-trans.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:
.lib "C:\ProgramFiles\Orcad\Capture\Library\PSpice\nom.lib" 
.inc "C:\ProgramFiles\Orcad\Capture\Library\PSpice\nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 50us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rectifier-SCHEMATIC1.net" 


.END
