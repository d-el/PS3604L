* D:\Radio\Devices\PS3608L\OrCad\CulerReg2.sch

* Schematics Version 9.2
* Tue Aug 09 01:20:36 2016



** Analysis setup **
.tran 20ns 30ms


* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "CulerReg2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
