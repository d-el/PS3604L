** Profile: "SCHEMATIC1-Bias"  [ D:\Radio\Devices\PS3608L\OrCad\reg-schematic1-bias.sim ] 

** Creating circuit file "reg-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OP
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\reg-SCHEMATIC1.net" 


.END
