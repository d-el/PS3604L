** Profile: "SCHEMATIC1-simpro"  [ d:\radio\devices\ps3608l\orcad\reg-schematic1-simpro.sim ] 

** Creating circuit file "reg-schematic1-simpro.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\programfiles\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10000ns 0 .001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\reg-SCHEMATIC1.net" 


.END
